`ifndef _constants_vh_
`define _constants_vh_

`define MIPS_CONTROL_ALU_B_SOURCE__IMMEDIATE 2'b00
`define MIPS_CONTROL_ALU_B_SOURCE__REGISTER_OUTPUT_2 2'b01
`define MIPS_CONTROL_ALU_B_SOURCE__SHIFT_IMMEDIATE 2'b10

`endif // _constants_vh_
